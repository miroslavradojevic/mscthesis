<?xml version="1.0" encoding="UTF-8" standalone="no"?>
<!-- Created with Inkscape (http://www.inkscape.org/) -->

<svg
   xmlns:dc="http://purl.org/dc/elements/1.1/"
   xmlns:cc="http://creativecommons.org/ns#"
   xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"
   xmlns:svg="http://www.w3.org/2000/svg"
   xmlns="http://www.w3.org/2000/svg"
   xmlns:sodipodi="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd"
   xmlns:inkscape="http://www.inkscape.org/namespaces/inkscape"
   width="744.09448819"
   height="1052.3622047"
   id="svg3797"
   version="1.1"
   inkscape:version="0.47 r22583"
   sodipodi:docname="auv-model.svg">
  <defs
     id="defs3799">
    <inkscape:perspective
       sodipodi:type="inkscape:persp3d"
       inkscape:vp_x="0 : 526.18109 : 1"
       inkscape:vp_y="0 : 1000 : 0"
       inkscape:vp_z="744.09448 : 526.18109 : 1"
       inkscape:persp3d-origin="372.04724 : 350.78739 : 1"
       id="perspective3805" />
    <inkscape:perspective
       id="perspective3732"
       inkscape:persp3d-origin="0.5 : 0.33333333 : 1"
       inkscape:vp_z="1 : 0.5 : 1"
       inkscape:vp_y="0 : 1000 : 0"
       inkscape:vp_x="0 : 0.5 : 1"
       sodipodi:type="inkscape:persp3d" />
    <marker
       inkscape:stockid="Arrow1Lstart"
       orient="auto"
       refY="0"
       refX="0"
       id="Arrow1Lstart"
       style="overflow:visible">
      <path
         id="path16098"
         d="M 0,0 5,-5 -12.5,0 5,5 0,0 z"
         style="fill-rule:evenodd;stroke:#000000;stroke-width:1pt;marker-start:none"
         transform="matrix(0.8,0,0,0.8,10,0)" />
    </marker>
    <marker
       inkscape:stockid="Arrow1Lend"
       orient="auto"
       refY="0"
       refX="0"
       id="Arrow1Lend"
       style="overflow:visible">
      <path
         id="path16101"
         d="M 0,0 5,-5 -12.5,0 5,5 0,0 z"
         style="fill-rule:evenodd;stroke:#000000;stroke-width:1pt;marker-start:none"
         transform="matrix(-0.8,0,0,-0.8,-10,0)" />
    </marker>
    <marker
       inkscape:stockid="Arrow1Mend"
       orient="auto"
       refY="0"
       refX="0"
       id="Arrow1Mend"
       style="overflow:visible">
      <path
         id="path16107"
         d="M 0,0 5,-5 -12.5,0 5,5 0,0 z"
         style="fill-rule:evenodd;stroke:#000000;stroke-width:1pt;marker-start:none"
         transform="matrix(-0.4,0,0,-0.4,-4,0)" />
    </marker>
    <marker
       inkscape:stockid="Arrow1Lstart"
       orient="auto"
       refY="0"
       refX="0"
       id="marker3742"
       style="overflow:visible">
      <path
         id="path3744"
         d="M 0,0 5,-5 -12.5,0 5,5 0,0 z"
         style="fill-rule:evenodd;stroke:#000000;stroke-width:1pt;marker-start:none"
         transform="matrix(0.8,0,0,0.8,10,0)" />
    </marker>
  </defs>
  <sodipodi:namedview
     id="base"
     pagecolor="#ffffff"
     bordercolor="#ffffff"
     borderopacity="0.0"
     inkscape:pageopacity="0.0"
     inkscape:pageshadow="0"
     inkscape:zoom="0.35"
     inkscape:cx="350"
     inkscape:cy="520"
     inkscape:document-units="px"
     inkscape:current-layer="layer1"
     showgrid="false"
     inkscape:window-width="1366"
     inkscape:window-height="693"
     inkscape:window-x="0"
     inkscape:window-y="24"
     inkscape:window-maximized="1" />
  <metadata
     id="metadata3802">
    <rdf:RDF>
      <cc:Work
         rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type
           rdf:resource="http://purl.org/dc/dcmitype/StillImage" />
        <dc:title></dc:title>
      </cc:Work>
    </rdf:RDF>
  </metadata>
  <g
     inkscape:label="Layer 1"
     inkscape:groupmode="layer"
     id="layer1">
    <path
       d="m -243.76073,1093.8806 0,-588.75706 1416.13193,0"
       style="fill:none;stroke:#231f20;stroke-width:9.87509918;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:22.92560005;stroke-opacity:1;stroke-dasharray:none"
       id="path13958-6" />
    <path
       d="m 1147.2979,532.60253 54.6067,-30.05064 -54.6067,-30.05639 0,60.10703"
       style="fill:#231f20;fill-opacity:1;fill-rule:evenodd;stroke:none"
       id="path13960-2" />
    <path
       d="m 344.10387,55.141886 59.84674,-17.37965 -17.3707,59.87767 -42.47604,-42.49802"
       style="fill:#231f20;fill-opacity:1;fill-rule:evenodd;stroke:none"
       id="path13962-5" />
    <path
       d="m -246.17693,546.17239 c 22.4805,0 40.7095,-18.24422 40.7095,-40.73622 0,-22.492 -18.229,-40.73044 -40.7095,-40.73044 -22.4861,0 -40.7151,18.23844 -40.7151,40.73044 0,22.492 18.229,40.73622 40.7151,40.73622 z"
       style="fill:none;stroke:#231f20;stroke-width:6.50721073;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:22.92560005;stroke-opacity:1;stroke-dasharray:none"
       id="path13964-4" />
    <path
       d="M -245.16633,499.93757 365.77987,73.731556"
       style="fill:none;stroke:#231f20;stroke-width:5.99866247;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:22.92560005;stroke-opacity:1;stroke-dasharray:none"
       id="path13970-4" />
    <g
       id="g15161-9"
       transform="matrix(0.26227731,-5.3927017,-5.1100985,-0.29800329,4085.2755,164.14279)"
       inkscape:transform-center-x="32.023884"
       inkscape:transform-center-y="31.397683">
      <path
         id="path13950-9"
         style="fill:#fff200;fill-opacity:1;fill-rule:evenodd;stroke:none"
         d="m -111.11535,690.69897 c -0.75479,-0.47824 -1.51283,-0.91745 -2.30341,-1.33063 -0.4815,-0.25377 -1.65923,-0.0182 -2.44655,0.28629 -7.6715,2.97361 -16.95018,12.7468 -20.96161,19.6928 -11.54955,20.00512 -20.81522,36.16472 -27.21139,48.87573 -4.58403,9.11601 -7.72356,19.78389 -9.65607,30.11342 l 3.5039,2.02361 3.50065,2.02035 c 7.98383,-6.83863 15.65208,-14.89078 21.25117,-23.41792 7.8114,-11.89441 17.17467,-27.99871 28.72422,-48.00058 4.00818,-6.94925 7.83417,-19.87498 6.57185,-28.00196 -0.12675,-0.83612 -0.51403,-1.97155 -0.97276,-2.26111" />
      <path
         id="path13952-3"
         style="fill:none;stroke:#231f20;stroke-width:0.39785165;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:22.92560005;stroke-opacity:1;stroke-dasharray:none"
         d="m -111.11535,690.69897 c -0.75479,-0.47824 -1.51283,-0.91745 -2.30341,-1.33063 -0.4815,-0.25377 -1.65923,-0.0182 -2.44655,0.28629 -7.6715,2.97361 -16.95018,12.7468 -20.96161,19.6928 -11.54955,20.00512 -20.81522,36.16472 -27.21139,48.87573 -4.58403,9.11601 -7.72356,19.78389 -9.65607,30.11342 l 3.5039,2.02361 3.50065,2.02035 c 7.98383,-6.83863 15.65208,-14.89078 21.25117,-23.41792 7.8114,-11.89441 17.17467,-27.99871 28.72422,-48.00058 4.00818,-6.94925 7.83417,-19.87498 6.57185,-28.00196 -0.12675,-0.83612 -0.51403,-1.97155 -0.97276,-2.26111 z" />
      <path
         id="path13954-6"
         style="fill:#0994dc;fill-opacity:1;fill-rule:evenodd;stroke:none"
         d="m -175.87741,787.20439 11.96924,6.91347 c 1.0541,0.60513 1.55837,1.71779 1.12242,2.46932 l -2.46282,4.26846 c -0.43596,0.75153 -1.64947,0.8719 -2.70032,0.26352 l -11.96923,-6.91021 c -1.05085,-0.60838 -1.55838,-1.71779 -1.12243,-2.47258 l 2.46282,-4.2652 c 0.43596,-0.75478 1.64947,-0.87191 2.70032,-0.26678" />
      <path
         id="path13956-0"
         style="fill:none;stroke:#231f20;stroke-width:0.39785165;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:22.92560005;stroke-opacity:1;stroke-dasharray:none"
         d="m -175.87741,787.20439 11.96924,6.91347 c 1.0541,0.60513 1.55837,1.71779 1.12242,2.46932 l -2.46282,4.26846 c -0.43596,0.75153 -1.64947,0.8719 -2.70032,0.26352 l -11.96923,-6.91021 c -1.05085,-0.60838 -1.55838,-1.71779 -1.12243,-2.47258 l 2.46282,-4.2652 c 0.43596,-0.75478 1.64947,-0.87191 2.70032,-0.26678 z" />
      <path
         id="path13980-5"
         style="fill:none;stroke:#231f20;stroke-width:0.92100805;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:22.92560005;stroke-opacity:1;stroke-dasharray:none"
         d="m -134.504,741.56253 c 1.54536,-2.67754 0.6279,-6.10662 -2.05289,-7.65198 -2.67755,-1.54861 -6.10662,-0.63116 -7.65524,2.04964 -1.54536,2.6808 -0.6279,6.10662 2.05289,7.65523 2.6808,1.54537 6.10662,0.62791 7.65524,-2.05289 z" />
      <path
         id="path13982-0"
         style="fill:#231f20;fill-opacity:1;fill-rule:evenodd;stroke:none"
         d="m -138.69437,739.26238 c 0.30907,-0.53681 0.12363,-1.22002 -0.40993,-1.53234 -0.53681,-0.30908 -1.22328,-0.12363 -1.53235,0.40992 -0.30907,0.53681 -0.12363,1.22328 0.40993,1.53235 0.53681,0.30907 1.22328,0.12363 1.53235,-0.40993" />
      <path
         id="path13984-2"
         style="fill:none;stroke:#231f20;stroke-width:0.92100805;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:22.92560005;stroke-opacity:1;stroke-dasharray:none"
         d="m -138.69437,739.26238 c 0.30907,-0.53681 0.12363,-1.22002 -0.40993,-1.53234 -0.53681,-0.30908 -1.22328,-0.12363 -1.53235,0.40992 -0.30907,0.53681 -0.12363,1.22328 0.40993,1.53235 0.53681,0.30907 1.22328,0.12363 1.53235,-0.40993 z" />
    </g>
    <path
       d="m -279.76433,1069.8141 30.035,54.635 30.0409,-54.635 -60.0759,0"
       style="fill:#231f20;fill-opacity:1;fill-rule:evenodd;stroke:none"
       id="path13960-4-9" />
    <path
       d="m -246.12303,232.74575 0,220.29295"
       style="fill:none;stroke:#231f20;stroke-width:1.39495432;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:22.92560005;stroke-opacity:1;stroke-dasharray:6.97477193, 4.18486316;stroke-dashoffset:0;marker-start:url(#Arrow1Lstart);marker-end:none"
       id="path13986-9-4" />
    <path
       d="m 274.40347,257.28021 0,435.64076"
       style="fill:none;stroke:#231f20;stroke-width:1.96166098;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:22.92560005;stroke-opacity:1;stroke-dasharray:9.80830537, 5.88498322;stroke-dashoffset:0"
       id="path13986-9-5-3" />
    <path
       d="M 271.58607,702.7784 858.73671,386.63041"
       style="fill:none;stroke:#231f20;stroke-width:2.86767602;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:22.92560005;stroke-opacity:1;stroke-dasharray:14.33838184, 8.60302911;stroke-dashoffset:0"
       id="path13986-9-5-5-5"
       sodipodi:nodetypes="cc" />
    <path
       d="M 269.86217,702.71851 1042.4072,450.94003"
       style="fill:none;stroke:#231f20;stroke-width:2.9354949;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:22.92560005;stroke-opacity:1;stroke-dasharray:14.6774763, 8.8064858;stroke-dashoffset:0"
       id="path13986-9-5-5-6-1"
       sodipodi:nodetypes="cc" />
    <g
       id="g15129-5"
       transform="matrix(1.765863,0,0,1.7667761,692.08631,-134.73814)">
      <path
         sodipodi:nodetypes="cc"
         id="path13990-1"
         style="fill:none;stroke:#231f20;stroke-width:0.97261995;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:22.92560005;stroke-opacity:1;stroke-dasharray:none"
         d="m -196.67938,237.44588 c 114.360227,19.39563 -0.35305,77.0244 -99.68862,68.09087" />
      <path
         id="path13960-6-6"
         style="fill:#231f20;fill-opacity:1;fill-rule:evenodd;stroke:none"
         d="m -291.6246,289.85923 -30.92351,17.00874 30.92351,17.01199 0,-34.02073" />
    </g>
    <path
       style="fill:none;stroke:#000000;stroke-width:3.20670176;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker-start:none;marker-end:url(#Arrow1Mend)"
       d="m 934.52931,480.40496 c 140.00439,-111.32276 -50.0017,-97.7468 -50.0017,-97.7468"
       id="path15321" />
    <text
       xml:space="preserve"
       style="font-size:86.79489899px;font-style:normal;font-weight:normal;fill:#000000;fill-opacity:1;stroke:none;font-family:Bitstream Vera Sans"
       x="248.98761"
       y="-6.4811492"
       id="text17397-7"
       transform="scale(0.99974156,1.0002585)"><tspan
         sodipodi:role="line"
         id="tspan17399-4"
         x="248.98761"
         y="-6.4811492"
         style="font-size:90px;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-family:BKM-cmr12;-inkscape-font-specification:BKM-cmr12">x (north)</tspan></text>
    <text
       xml:space="preserve"
       style="font-size:70.65277863px;font-style:normal;font-weight:normal;fill:#000000;fill-opacity:1;stroke:none;font-family:Bitstream Vera Sans"
       x="994.62659"
       y="598.34674"
       id="text17397-6-3"
       transform="scale(0.99974156,1.0002585)"><tspan
         sodipodi:role="line"
         id="tspan17399-9-1"
         x="994.62659"
         y="598.34674"
         style="font-size:90px;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-family:BKM-cmr12;-inkscape-font-specification:BKM-cmr12">x (east)</tspan></text>
    <text
       xml:space="preserve"
       style="font-size:70.65277863px;font-style:normal;font-weight:normal;fill:#000000;fill-opacity:1;stroke:none;font-family:Bitstream Vera Sans"
       x="-205.03265"
       y="988.69611"
       id="text17397-8-4"
       transform="scale(0.99974156,1.0002585)"><tspan
         sodipodi:role="line"
         id="tspan17399-3-6"
         x="-205.03265"
         y="988.69611"
         style="font-size:90px;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-family:BKM-cmr12;-inkscape-font-specification:BKM-cmr12">z (depth)</tspan></text>
    <text
       xml:space="preserve"
       style="font-size:70.65277863px;font-style:normal;font-weight:normal;fill:#000000;fill-opacity:1;stroke:none;font-family:Bitstream Vera Sans"
       x="361.55756"
       y="249.28941"
       id="text17397-6-8"
       transform="scale(0.99974156,1.0002585)"><tspan
         sodipodi:role="line"
         id="tspan17399-9-3"
         x="361.55756"
         y="249.28941"
         style="font-size:90px;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-family:BKM-cmr12;-inkscape-font-specification:BKM-cmr12"> (yaw)</tspan></text>
    <text
       xml:space="preserve"
       style="font-size:70.65277863px;font-style:normal;font-weight:normal;fill:#000000;fill-opacity:1;stroke:none;font-family:Bitstream Vera Sans"
       x="1038.0211"
       y="380.50168"
       id="text17397-6-8-5"
       transform="scale(0.99974156,1.0002585)"><tspan
         sodipodi:role="line"
         id="tspan17399-9-3-0"
         x="1038.0211"
         y="380.50168"
         style="font-size:90px;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-family:BKM-cmr12;-inkscape-font-specification:BKM-cmr12"> (pitch)</tspan></text>
    <text
       xml:space="preserve"
       style="font-size:94.05136871px;font-style:normal;font-weight:normal;fill:#000000;fill-opacity:1;stroke:none;font-family:Bitstream Vera Sans"
       x="317.13275"
       y="242.52599"
       id="text19778"
       transform="scale(0.99974156,1.0002585)"><tspan
         sodipodi:role="line"
         id="tspan19780"
         x="317.13275"
         y="242.52599">ψ</tspan></text>
    <text
       style="font-size:88.28483582px"
       y="393.35797"
       x="1006.8054"
       id="text19648"
       transform="scale(0.99974156,1.0002585)">
      <tspan
         style="font-size:87.95523834px;font-variant:normal;font-weight:normal;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;font-family:CMMI12;-inkscape-font-specification:CMMI12"
         x="1006.8054"
         y="393.35797"
         id="tspan19650">θ</tspan>
    </text>
    <path
       d="m 562.64681,705.78754 0,366.68856"
       style="fill:none;stroke:#231f20;stroke-width:2.31787658;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:22.92560005;stroke-opacity:1;stroke-dasharray:11.58938302, 6.95362981;stroke-dashoffset:0;marker-start:url(#Arrow1Lstart);marker-end:url(#Arrow1Lend)"
       id="path13986-9-3" />
    <text
       xml:space="preserve"
       style="font-size:70.65277863px;font-style:normal;font-weight:normal;fill:#000000;fill-opacity:1;stroke:none;font-family:Bitstream Vera Sans"
       x="615.16077"
       y="745.80847"
       id="text17397-8-8"
       transform="scale(0.99974156,1.0002585)"><tspan
         sodipodi:role="line"
         id="tspan17399-3-1"
         x="615.16077"
         y="745.80847"
         style="font-size:90px;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-family:BKM-cmr12;-inkscape-font-specification:BKM-cmr12">a (altitude)</tspan></text>
    <path
       style="fill:#000000;fill-opacity:1;stroke:#000000;stroke-width:2.58362532;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0"
       id="path21308-9"
       d="m -169.59023,1113.5774 c 15.6032,-2.6936 30.6573,-7.0906 45.5545,-11.4221 25.054901,-8.5202 51.536601,-14.2784 76.958801,-22.0806 32.6549,-11.8655 65.5639,-23.3367 98.1234,-35.3472 20.0684,-8.1547 41.8113,-13.5803 62.573299,-20.5694 10.7662,-3.9256 22.2967,-6.2997 34.2289,-6.9939 14.1226,-0.5014 28.2805,-0.2678 42.4157,-0.1976 15.6385,-0.035 31.2772,0.041 46.9155,0.012 16.3408,-0.794 32.3345,1.5399 48.4433,3.0854 18.7863,2.2944 37.1806,6.2999 55.5037,10.1198 17.7803,2.9322 34.9459,7.5246 52.21904,11.7582 18.0583,3.9422 36.2254,7.554 54.2811,11.5058 15.9123,3.2439 31.989,6.0383 47.8799,9.3349 14.7087,3.7666 29.5024,7.3123 44.7024,9.8206 2.4472,0.4435 4.9244,0.8036 7.3415,1.3299 5.0943,1.1088 10.0247,2.5993 15.0854,3.7895 6.8573,1.6129 13.8661,2.7567 20.8041,4.1548 13.671,2.3231 27.201,5.0818 40.98,7.051 12.7893,3.1071 25.6375,6.0002 38.5796,8.7298 14.7155,3.1643 29.9183,4.3717 44.9717,6.2155 12.5176,2.3354 25.1119,4.1884 37.9661,5.0647 11.4597,0.5977 22.958,0.6283 34.441,0.6245 12.3838,0.018 24.7674,0.021 37.151,-0.044 10.8808,0.044 21.7616,-0.039 32.6421,-0.09 8.6424,0.2816 17.1002,-0.1679 25.6556,-0.9073 11.7012,-0.4357 23.046,-2.5106 34.5082,-4.0941 14.6865,-2.5062 29.0659,-5.8744 43.5102,-9.041 15.0489,-2.71 29.9179,-5.8929 44.789,-9.0865 14.74349,-3.6215 29.93129,-5.6987 45.11169,-7.9383 13.8755,-1.8698 27.9528,-2.5761 42.0176,-3.0908 10.1083,-0.2657 20.2222,-0.27 30.335,-0.2666 5.949,0 3.0069,0 8.8262,0 0,0 -42.4322,22.8412 -42.4322,22.8412 l 0,0 c -5.7645,-0.023 -2.8494,-0.018 -8.7455,-0.032 -9.9762,-0.018 -19.9579,-0.023 -29.9275,0.2771 -13.8571,0.4674 -27.7014,1.327 -41.315,3.3941 -15.03609,2.1074 -29.88929,4.6768 -44.52239,8.0332 -14.9471,3.1811 -29.8625,6.4197 -44.9526,9.2151 -14.5786,3.2087 -29.1341,6.5489 -44.0253,8.8862 -11.6059,1.8035 -23.2628,3.2816 -35.0888,4.0426 -8.6849,0.7736 -17.3938,0.6818 -26.132,0.6005 -10.7849,-0.046 -21.5703,-0.1254 -32.3554,-0.06 -12.3836,-0.041 -24.7665,0.023 -37.1501,0.021 -11.6055,-0.064 -23.2353,-0.026 -34.7929,-0.9318 -12.7648,-1.172 -25.1926,-3.3764 -37.739,-5.4319 -15.2637,-1.7903 -30.5773,-3.4322 -45.5132,-6.4645 -12.862,-2.6348 -25.4187,-5.9916 -38.3148,-8.5294 -13.7919,-2.203 -27.4617,-4.8064 -41.1751,-7.2585 -14.3884,-2.9431 -28.4962,-6.5137 -42.9521,-9.2522 -15.1603,-2.8073 -30.0188,-6.3661 -44.8891,-9.9095 -15.8183,-3.2497 -31.7053,-6.3145 -47.5098,-9.6025 -18.051,-4.0022 -36.32994,-7.4052 -54.29694,-11.6188 -17.3062,-4.1261 -34.5132,-8.5367 -52.2519,-11.5586 -18.1258,-3.8139 -36.3084,-7.9155 -55.0467,-9.666 -16.0899,-1.4879 -32.1108,-3.2597 -48.3921,-2.5261 -15.5571,-0.06 -31.1148,-0.044 -46.6719,-0.1434 -14.2511,0.042 -28.5503,-0.093 -42.7493,0.9367 -11.404599,1.3103 -22.333399,3.8276 -32.743299,7.5734 -20.3654,6.2635 -41.0341,12.0259 -60.5981,19.6433 -32.7126,11.9475 -65.6795,23.5128 -98.5283,35.2488 -25.904701,7.7314 -52.523501,14.1051 -78.019001,22.6165 -15.621,4.4484 -31.2724,8.9305 -47.4779,12.0839 0,0 41.7927,-23.852 41.7927,-23.852 z" />
    <path
       d="m -619.89783,503.32355 c 36.9041,46.42131 38.4349,-40.31271 73.3813,0 36.8718,46.26261 37.7466,-40.47145 72.693,0 36.872,46.26261 38.0773,-40.47145 73.0186,0 36.8776,46.26261 38.0775,-40.47145 73.0239,0 36.8718,46.26261 38.0775,-40.47145 73.0238,0"
       style="fill:none;stroke:#00adef;stroke-width:5.7605114;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:22.92560005;stroke-opacity:1;stroke-dasharray:none"
       id="path21709-4" />
  </g>
</svg>
